module file_reg_top (       
);

        

endmodule
