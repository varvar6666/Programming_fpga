module part_2_top_module ();

// write code here


endmodule