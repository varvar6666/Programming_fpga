module part_5_top_module (input [31:0]a, input [31:0]b, input sub, output [31:0] sum);

    // write code here

endmodule