module ram_top(
);
    

endmodule
