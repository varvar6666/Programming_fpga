module part_4_top_module (input [31:0]a, input [31:0]b, input cin, output [31:0] sum, output cout);

    // write code here

endmodule