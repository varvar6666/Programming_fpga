module lut_top (

);
    

endmodule
