module sevenseg_top(
);
    

endmodule
