module sync_top(
);
    

endmodule
