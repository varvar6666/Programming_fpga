module part_1_top_module (input clk, input d, output q );

    // write code here


endmodule