module m_not (input wire in, output wire out);
assign out = ~in;
endmodule