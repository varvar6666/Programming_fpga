module part_1_top_module ();

// write code here


endmodule