module part_3_top_module ();

// write code here


endmodule