module part_5_top_module ();

// write code here

endmodule