module rom_top(
);
    

endmodule
