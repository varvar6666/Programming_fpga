module part_4_top_module ();

// write code here


endmodule