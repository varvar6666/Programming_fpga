`define MODULE_NAME Integer_Multiplier_Top
`define UNSIGNED_A
`define UNSIGNED_B
`define DATA_B
`define LUT
`define NON_PIPELINE
