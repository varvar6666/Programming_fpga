
module part_2_top_module (input [7:0]d, input [1:0]sel, input clk, output reg [7:0]q);

    // write code here

endmodule