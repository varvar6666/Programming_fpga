// Часть 1: Комбинационная схема
// Анализируя временную диаграмму, это выглядит как логическая функция
module part1_combinational(
    input a,
    input b,
    input c,
    output y
);

// Логика на основе анализа временной диаграммы
assign y = c;

endmodule
