parameter WIDTH_B = 8;
parameter WIDTH_A = 8;
